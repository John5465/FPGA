module Test_Led(
	CLK,RSTn,
	led
);

input CLK;
input RSTn;
output led;

assign led = 1'b1;	


endmodule