module Speed_Select();

endmodule