module Uart_Tx();

endmodule