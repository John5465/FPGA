module B(a,b,y); //两个数相乘的模块
input [1:0]a;
input [1:0]b;
output [3:0]y;
assign y=a*b ;
endmodule 