module top_calc(
clk,rst_n,
y
);

input clk;
input rst_n;
output y;


endmodule